interface intf;
  
  logic reset;
  logic clk;
  logic d;
  logic q;
  logic qbar;
  
endinterface
